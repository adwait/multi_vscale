//A 4-core system!
`define NUM_CORES 2
`define CORE_IDX_WIDTH 1
